module sub_module #(
  /*AUTOINOUTPARAM*/
)(
  /*AUTOARG*/
);

  /*AUTOVARIABLE*/

  /*AUTOINST*/

endmodule
